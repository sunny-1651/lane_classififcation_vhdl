LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.HDLLaneDetector_pkg.ALL;

ENTITY Horizontal_Padder IS
  PORT( clk                               :   IN    std_logic;
        reset                             :   IN    std_logic;
        enb                               :   IN    std_logic;
        dataVectorIn                      :   IN    vector_of_std_logic_vector8(0 TO 15);  -- uint8 [16]
        horPadCount                       :   IN    std_logic_vector(10 DOWNTO 0);  -- ufix11
        padShift                          :   IN    std_logic;
        dataVector                        :   OUT   vector_of_std_logic_vector8(0 TO 15)  -- uint8 [16]
        );
END Horizontal_Padder;


ARCHITECTURE rtl OF Horizontal_Padder IS

  -- Signals
  SIGNAL horPadCount_unsigned             : unsigned(10 DOWNTO 0);  -- ufix11
  SIGNAL dataVectorIn_unsigned            : vector_of_unsigned8(0 TO 15);  -- uint8 [16]
  SIGNAL DataMuxIn1                       : vector_of_unsigned8(0 TO 15);  -- uint8 [16]
  SIGNAL DataMuxIn1_0                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_1                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_2                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_3                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_4                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_5                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_6                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_7                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_8                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_9                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_10                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_11                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_12                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_13                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_14                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn1_15                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_1                   : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg                   : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_out_2                   : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_3                   : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_4                   : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_5                   : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_6                   : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_7                   : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_8                   : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_9                   : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_10                  : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_11                  : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_12                  : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_13                  : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_14                  : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_15                  : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_16                  : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_1                 : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_2                 : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_3                 : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_4                 : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_5                 : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_6                 : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_7                 : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_8                 : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_9                 : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_10                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_11                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_12                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_13                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_14                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_15                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL DataMuxIn1_16                    : vector_of_unsigned8(0 TO 15);  -- uint8 [16]
  SIGNAL intdelay_out_1_1                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_16                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_out_2_1                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_3_1                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_4_1                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_5_1                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_6_1                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_7_1                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_8_1                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_9_1                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_10_1                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_11_1                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_12_1                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_13_1                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_14_1                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_15_1                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_16_1                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_17                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_18                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_19                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_20                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_21                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_22                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_23                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_24                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_25                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_26                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_27                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_28                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_29                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_30                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_31                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL DataMuxIn2                       : vector_of_unsigned8(0 TO 15);  -- uint8 [16]
  SIGNAL DataMuxIn3                       : vector_of_unsigned8(0 TO 15);  -- uint8 [16]
  SIGNAL DataMuxIn4                       : vector_of_unsigned8(0 TO 15);  -- uint8 [16]
  SIGNAL DataMuxIn4_0                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_1                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_2                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_3                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_4                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_5                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_6                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_7                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_8                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_9                     : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_10                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_11                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_12                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_13                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_14                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL DataMuxIn4_15                    : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_1_2                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_32                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_out_2_2                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_3_2                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_4_2                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_5_2                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_6_2                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_7_2                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_8_2                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_9_2                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_10_2                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_11_2                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_12_2                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_13_2                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_14_2                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_15_2                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_16_2                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_33                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_34                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_35                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_36                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_37                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_38                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_39                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_40                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_41                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_42                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_43                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_44                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_45                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_46                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_47                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL DataMuxIn5                       : vector_of_unsigned8(0 TO 15);  -- uint8 [16]
  SIGNAL intdelay_out_1_3                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_48                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_out_2_3                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_3_3                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_4_3                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_5_3                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_6_3                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_7_3                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_8_3                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_9_3                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_10_3                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_11_3                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_12_3                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_13_3                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_14_3                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_15_3                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_16_3                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_49                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_50                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_51                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_52                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_53                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_54                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_55                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_56                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_57                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_58                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_59                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_60                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_61                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_62                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_63                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL DataMuxIn6                       : vector_of_unsigned8(0 TO 15);  -- uint8 [16]
  SIGNAL intdelay_out_1_4                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_64                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_out_2_4                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_3_4                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_4_4                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_5_4                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_6_4                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_7_4                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_8_4                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_9_4                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_10_4                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_11_4                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_12_4                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_13_4                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_14_4                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_15_4                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_16_4                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_65                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_66                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_67                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_68                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_69                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_70                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_71                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_72                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_73                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_74                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_75                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_76                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_77                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_78                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_79                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL DataMuxIn7                       : vector_of_unsigned8(0 TO 15);  -- uint8 [16]
  SIGNAL intdelay_out_1_5                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_80                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_out_2_5                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_3_5                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_4_5                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_5_5                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_6_5                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_7_5                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_8_5                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_9_5                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_10_5                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_11_5                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_12_5                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_13_5                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_14_5                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_15_5                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_16_5                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_81                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_82                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_83                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_84                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_85                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_86                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_87                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_88                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_89                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_90                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_91                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_92                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_93                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_94                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_95                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL DataMuxIn8                       : vector_of_unsigned8(0 TO 15);  -- uint8 [16]
  SIGNAL intdelay_out_1_6                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_96                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_out_2_6                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_3_6                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_4_6                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_5_6                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_6_6                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_7_6                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_8_6                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_9_6                 : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_10_6                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_11_6                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_12_6                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_13_6                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_14_6                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_15_6                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_out_16_6                : unsigned(7 DOWNTO 0);  -- uint8
  SIGNAL intdelay_1_reg_97                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_98                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_99                : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_100               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_101               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_102               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_103               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_104               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_105               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_106               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_107               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_108               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_109               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_110               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL intdelay_1_reg_111               : vector_of_unsigned8(0 TO 1);  -- ufix8 [2]
  SIGNAL DataMuxIn9                       : vector_of_unsigned8(0 TO 15);  -- uint8 [16]
  SIGNAL dataVector_tmp                   : vector_of_unsigned8(0 TO 15);  -- uint8 [16]

BEGIN
  horPadCount_unsigned <= unsigned(horPadCount);

  outputgen1: FOR k IN 0 TO 15 GENERATE
    dataVectorIn_unsigned(k) <= unsigned(dataVectorIn(k));
  END GENERATE;

  reg_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        DataMuxIn1 <= (OTHERS => to_unsigned(16#00#, 8));
      ELSIF enb = '1' AND padShift = '1' THEN
        DataMuxIn1 <= dataVectorIn_unsigned;
      END IF;
    END IF;
  END PROCESS reg_process;


  DataMuxIn1_0 <= DataMuxIn1(0);

  intdelay_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        intdelay_1_reg <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_1 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_2 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_3 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_4 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_5 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_6 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_7 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_8 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_9 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_10 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_11 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_12 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_13 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_14 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_15 <= (OTHERS => to_unsigned(16#00#, 8));
      ELSIF enb = '1' AND padShift = '1' THEN
        intdelay_1_reg(0) <= DataMuxIn1_0;
        intdelay_1_reg(1) <= intdelay_1_reg(0);
        intdelay_1_reg_1(0) <= DataMuxIn1_1;
        intdelay_1_reg_1(1) <= intdelay_1_reg_1(0);
        intdelay_1_reg_2(0) <= DataMuxIn1_2;
        intdelay_1_reg_2(1) <= intdelay_1_reg_2(0);
        intdelay_1_reg_3(0) <= DataMuxIn1_3;
        intdelay_1_reg_3(1) <= intdelay_1_reg_3(0);
        intdelay_1_reg_4(0) <= DataMuxIn1_4;
        intdelay_1_reg_4(1) <= intdelay_1_reg_4(0);
        intdelay_1_reg_5(0) <= DataMuxIn1_5;
        intdelay_1_reg_5(1) <= intdelay_1_reg_5(0);
        intdelay_1_reg_6(0) <= DataMuxIn1_6;
        intdelay_1_reg_6(1) <= intdelay_1_reg_6(0);
        intdelay_1_reg_7(0) <= DataMuxIn1_7;
        intdelay_1_reg_7(1) <= intdelay_1_reg_7(0);
        intdelay_1_reg_8(0) <= DataMuxIn1_8;
        intdelay_1_reg_8(1) <= intdelay_1_reg_8(0);
        intdelay_1_reg_9(0) <= DataMuxIn1_9;
        intdelay_1_reg_9(1) <= intdelay_1_reg_9(0);
        intdelay_1_reg_10(0) <= DataMuxIn1_10;
        intdelay_1_reg_10(1) <= intdelay_1_reg_10(0);
        intdelay_1_reg_11(0) <= DataMuxIn1_11;
        intdelay_1_reg_11(1) <= intdelay_1_reg_11(0);
        intdelay_1_reg_12(0) <= DataMuxIn1_12;
        intdelay_1_reg_12(1) <= intdelay_1_reg_12(0);
        intdelay_1_reg_13(0) <= DataMuxIn1_13;
        intdelay_1_reg_13(1) <= intdelay_1_reg_13(0);
        intdelay_1_reg_14(0) <= DataMuxIn1_14;
        intdelay_1_reg_14(1) <= intdelay_1_reg_14(0);
        intdelay_1_reg_15(0) <= DataMuxIn1_15;
        intdelay_1_reg_15(1) <= intdelay_1_reg_15(0);
      END IF;
    END IF;
  END PROCESS intdelay_1_process;

  intdelay_out_1 <= intdelay_1_reg(1);
  intdelay_out_2 <= intdelay_1_reg_1(1);
  intdelay_out_3 <= intdelay_1_reg_2(1);
  intdelay_out_4 <= intdelay_1_reg_3(1);
  intdelay_out_5 <= intdelay_1_reg_4(1);
  intdelay_out_6 <= intdelay_1_reg_5(1);
  intdelay_out_7 <= intdelay_1_reg_6(1);
  intdelay_out_8 <= intdelay_1_reg_7(1);
  intdelay_out_9 <= intdelay_1_reg_8(1);
  intdelay_out_10 <= intdelay_1_reg_9(1);
  intdelay_out_11 <= intdelay_1_reg_10(1);
  intdelay_out_12 <= intdelay_1_reg_11(1);
  intdelay_out_13 <= intdelay_1_reg_12(1);
  intdelay_out_14 <= intdelay_1_reg_13(1);
  intdelay_out_15 <= intdelay_1_reg_14(1);
  intdelay_out_16 <= intdelay_1_reg_15(1);

  DataMuxIn1_1 <= DataMuxIn1(1);

  DataMuxIn1_2 <= DataMuxIn1(2);

  DataMuxIn1_3 <= DataMuxIn1(3);

  DataMuxIn1_4 <= DataMuxIn1(4);

  DataMuxIn1_5 <= DataMuxIn1(5);

  DataMuxIn1_6 <= DataMuxIn1(6);

  DataMuxIn1_7 <= DataMuxIn1(7);

  DataMuxIn1_8 <= DataMuxIn1(8);

  DataMuxIn1_9 <= DataMuxIn1(9);

  DataMuxIn1_10 <= DataMuxIn1(10);

  DataMuxIn1_11 <= DataMuxIn1(11);

  DataMuxIn1_12 <= DataMuxIn1(12);

  DataMuxIn1_13 <= DataMuxIn1(13);

  DataMuxIn1_14 <= DataMuxIn1(14);

  DataMuxIn1_15 <= DataMuxIn1(15);

  DataMuxIn1_16(0) <= intdelay_out_1;
  DataMuxIn1_16(1) <= intdelay_out_2;
  DataMuxIn1_16(2) <= intdelay_out_3;
  DataMuxIn1_16(3) <= intdelay_out_4;
  DataMuxIn1_16(4) <= intdelay_out_5;
  DataMuxIn1_16(5) <= intdelay_out_6;
  DataMuxIn1_16(6) <= intdelay_out_7;
  DataMuxIn1_16(7) <= intdelay_out_8;
  DataMuxIn1_16(8) <= intdelay_out_9;
  DataMuxIn1_16(9) <= intdelay_out_10;
  DataMuxIn1_16(10) <= intdelay_out_11;
  DataMuxIn1_16(11) <= intdelay_out_12;
  DataMuxIn1_16(12) <= intdelay_out_13;
  DataMuxIn1_16(13) <= intdelay_out_14;
  DataMuxIn1_16(14) <= intdelay_out_15;
  DataMuxIn1_16(15) <= intdelay_out_16;

  intdelay_1_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        intdelay_1_reg_16 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_17 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_18 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_19 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_20 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_21 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_22 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_23 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_24 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_25 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_26 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_27 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_28 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_29 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_30 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_31 <= (OTHERS => to_unsigned(16#00#, 8));
      ELSIF enb = '1' AND padShift = '1' THEN
        intdelay_1_reg_16(0) <= intdelay_out_1;
        intdelay_1_reg_16(1) <= intdelay_1_reg_16(0);
        intdelay_1_reg_17(0) <= intdelay_out_2;
        intdelay_1_reg_17(1) <= intdelay_1_reg_17(0);
        intdelay_1_reg_18(0) <= intdelay_out_3;
        intdelay_1_reg_18(1) <= intdelay_1_reg_18(0);
        intdelay_1_reg_19(0) <= intdelay_out_4;
        intdelay_1_reg_19(1) <= intdelay_1_reg_19(0);
        intdelay_1_reg_20(0) <= intdelay_out_5;
        intdelay_1_reg_20(1) <= intdelay_1_reg_20(0);
        intdelay_1_reg_21(0) <= intdelay_out_6;
        intdelay_1_reg_21(1) <= intdelay_1_reg_21(0);
        intdelay_1_reg_22(0) <= intdelay_out_7;
        intdelay_1_reg_22(1) <= intdelay_1_reg_22(0);
        intdelay_1_reg_23(0) <= intdelay_out_8;
        intdelay_1_reg_23(1) <= intdelay_1_reg_23(0);
        intdelay_1_reg_24(0) <= intdelay_out_9;
        intdelay_1_reg_24(1) <= intdelay_1_reg_24(0);
        intdelay_1_reg_25(0) <= intdelay_out_10;
        intdelay_1_reg_25(1) <= intdelay_1_reg_25(0);
        intdelay_1_reg_26(0) <= intdelay_out_11;
        intdelay_1_reg_26(1) <= intdelay_1_reg_26(0);
        intdelay_1_reg_27(0) <= intdelay_out_12;
        intdelay_1_reg_27(1) <= intdelay_1_reg_27(0);
        intdelay_1_reg_28(0) <= intdelay_out_13;
        intdelay_1_reg_28(1) <= intdelay_1_reg_28(0);
        intdelay_1_reg_29(0) <= intdelay_out_14;
        intdelay_1_reg_29(1) <= intdelay_1_reg_29(0);
        intdelay_1_reg_30(0) <= intdelay_out_15;
        intdelay_1_reg_30(1) <= intdelay_1_reg_30(0);
        intdelay_1_reg_31(0) <= intdelay_out_16;
        intdelay_1_reg_31(1) <= intdelay_1_reg_31(0);
      END IF;
    END IF;
  END PROCESS intdelay_1_1_process;

  intdelay_out_1_1 <= intdelay_1_reg_16(1);
  intdelay_out_2_1 <= intdelay_1_reg_17(1);
  intdelay_out_3_1 <= intdelay_1_reg_18(1);
  intdelay_out_4_1 <= intdelay_1_reg_19(1);
  intdelay_out_5_1 <= intdelay_1_reg_20(1);
  intdelay_out_6_1 <= intdelay_1_reg_21(1);
  intdelay_out_7_1 <= intdelay_1_reg_22(1);
  intdelay_out_8_1 <= intdelay_1_reg_23(1);
  intdelay_out_9_1 <= intdelay_1_reg_24(1);
  intdelay_out_10_1 <= intdelay_1_reg_25(1);
  intdelay_out_11_1 <= intdelay_1_reg_26(1);
  intdelay_out_12_1 <= intdelay_1_reg_27(1);
  intdelay_out_13_1 <= intdelay_1_reg_28(1);
  intdelay_out_14_1 <= intdelay_1_reg_29(1);
  intdelay_out_15_1 <= intdelay_1_reg_30(1);
  intdelay_out_16_1 <= intdelay_1_reg_31(1);

  DataMuxIn2(0) <= intdelay_out_1_1;
  DataMuxIn2(1) <= intdelay_out_2_1;
  DataMuxIn2(2) <= intdelay_out_3_1;
  DataMuxIn2(3) <= intdelay_out_4_1;
  DataMuxIn2(4) <= intdelay_out_5_1;
  DataMuxIn2(5) <= intdelay_out_6_1;
  DataMuxIn2(6) <= intdelay_out_7_1;
  DataMuxIn2(7) <= intdelay_out_8_1;
  DataMuxIn2(8) <= intdelay_out_9_1;
  DataMuxIn2(9) <= intdelay_out_10_1;
  DataMuxIn2(10) <= intdelay_out_11_1;
  DataMuxIn2(11) <= intdelay_out_12_1;
  DataMuxIn2(12) <= intdelay_out_13_1;
  DataMuxIn2(13) <= intdelay_out_14_1;
  DataMuxIn2(14) <= intdelay_out_15_1;
  DataMuxIn2(15) <= intdelay_out_16_1;

  reg_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        DataMuxIn3 <= (OTHERS => to_unsigned(16#00#, 8));
      ELSIF enb = '1' AND padShift = '1' THEN
        DataMuxIn3 <= DataMuxIn2;
      END IF;
    END IF;
  END PROCESS reg_1_process;


  reg_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        DataMuxIn4 <= (OTHERS => to_unsigned(16#00#, 8));
      ELSIF enb = '1' AND padShift = '1' THEN
        DataMuxIn4 <= DataMuxIn3;
      END IF;
    END IF;
  END PROCESS reg_2_process;


  DataMuxIn4_0 <= DataMuxIn4(0);

  intdelay_1_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        intdelay_1_reg_32 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_33 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_34 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_35 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_36 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_37 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_38 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_39 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_40 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_41 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_42 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_43 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_44 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_45 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_46 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_47 <= (OTHERS => to_unsigned(16#00#, 8));
      ELSIF enb = '1' AND padShift = '1' THEN
        intdelay_1_reg_32(0) <= DataMuxIn4_0;
        intdelay_1_reg_32(1) <= intdelay_1_reg_32(0);
        intdelay_1_reg_33(0) <= DataMuxIn4_1;
        intdelay_1_reg_33(1) <= intdelay_1_reg_33(0);
        intdelay_1_reg_34(0) <= DataMuxIn4_2;
        intdelay_1_reg_34(1) <= intdelay_1_reg_34(0);
        intdelay_1_reg_35(0) <= DataMuxIn4_3;
        intdelay_1_reg_35(1) <= intdelay_1_reg_35(0);
        intdelay_1_reg_36(0) <= DataMuxIn4_4;
        intdelay_1_reg_36(1) <= intdelay_1_reg_36(0);
        intdelay_1_reg_37(0) <= DataMuxIn4_5;
        intdelay_1_reg_37(1) <= intdelay_1_reg_37(0);
        intdelay_1_reg_38(0) <= DataMuxIn4_6;
        intdelay_1_reg_38(1) <= intdelay_1_reg_38(0);
        intdelay_1_reg_39(0) <= DataMuxIn4_7;
        intdelay_1_reg_39(1) <= intdelay_1_reg_39(0);
        intdelay_1_reg_40(0) <= DataMuxIn4_8;
        intdelay_1_reg_40(1) <= intdelay_1_reg_40(0);
        intdelay_1_reg_41(0) <= DataMuxIn4_9;
        intdelay_1_reg_41(1) <= intdelay_1_reg_41(0);
        intdelay_1_reg_42(0) <= DataMuxIn4_10;
        intdelay_1_reg_42(1) <= intdelay_1_reg_42(0);
        intdelay_1_reg_43(0) <= DataMuxIn4_11;
        intdelay_1_reg_43(1) <= intdelay_1_reg_43(0);
        intdelay_1_reg_44(0) <= DataMuxIn4_12;
        intdelay_1_reg_44(1) <= intdelay_1_reg_44(0);
        intdelay_1_reg_45(0) <= DataMuxIn4_13;
        intdelay_1_reg_45(1) <= intdelay_1_reg_45(0);
        intdelay_1_reg_46(0) <= DataMuxIn4_14;
        intdelay_1_reg_46(1) <= intdelay_1_reg_46(0);
        intdelay_1_reg_47(0) <= DataMuxIn4_15;
        intdelay_1_reg_47(1) <= intdelay_1_reg_47(0);
      END IF;
    END IF;
  END PROCESS intdelay_1_2_process;

  intdelay_out_1_2 <= intdelay_1_reg_32(1);
  intdelay_out_2_2 <= intdelay_1_reg_33(1);
  intdelay_out_3_2 <= intdelay_1_reg_34(1);
  intdelay_out_4_2 <= intdelay_1_reg_35(1);
  intdelay_out_5_2 <= intdelay_1_reg_36(1);
  intdelay_out_6_2 <= intdelay_1_reg_37(1);
  intdelay_out_7_2 <= intdelay_1_reg_38(1);
  intdelay_out_8_2 <= intdelay_1_reg_39(1);
  intdelay_out_9_2 <= intdelay_1_reg_40(1);
  intdelay_out_10_2 <= intdelay_1_reg_41(1);
  intdelay_out_11_2 <= intdelay_1_reg_42(1);
  intdelay_out_12_2 <= intdelay_1_reg_43(1);
  intdelay_out_13_2 <= intdelay_1_reg_44(1);
  intdelay_out_14_2 <= intdelay_1_reg_45(1);
  intdelay_out_15_2 <= intdelay_1_reg_46(1);
  intdelay_out_16_2 <= intdelay_1_reg_47(1);

  DataMuxIn4_1 <= DataMuxIn4(1);

  DataMuxIn4_2 <= DataMuxIn4(2);

  DataMuxIn4_3 <= DataMuxIn4(3);

  DataMuxIn4_4 <= DataMuxIn4(4);

  DataMuxIn4_5 <= DataMuxIn4(5);

  DataMuxIn4_6 <= DataMuxIn4(6);

  DataMuxIn4_7 <= DataMuxIn4(7);

  DataMuxIn4_8 <= DataMuxIn4(8);

  DataMuxIn4_9 <= DataMuxIn4(9);

  DataMuxIn4_10 <= DataMuxIn4(10);

  DataMuxIn4_11 <= DataMuxIn4(11);

  DataMuxIn4_12 <= DataMuxIn4(12);

  DataMuxIn4_13 <= DataMuxIn4(13);

  DataMuxIn4_14 <= DataMuxIn4(14);

  DataMuxIn4_15 <= DataMuxIn4(15);

  DataMuxIn5(0) <= intdelay_out_1_2;
  DataMuxIn5(1) <= intdelay_out_2_2;
  DataMuxIn5(2) <= intdelay_out_3_2;
  DataMuxIn5(3) <= intdelay_out_4_2;
  DataMuxIn5(4) <= intdelay_out_5_2;
  DataMuxIn5(5) <= intdelay_out_6_2;
  DataMuxIn5(6) <= intdelay_out_7_2;
  DataMuxIn5(7) <= intdelay_out_8_2;
  DataMuxIn5(8) <= intdelay_out_9_2;
  DataMuxIn5(9) <= intdelay_out_10_2;
  DataMuxIn5(10) <= intdelay_out_11_2;
  DataMuxIn5(11) <= intdelay_out_12_2;
  DataMuxIn5(12) <= intdelay_out_13_2;
  DataMuxIn5(13) <= intdelay_out_14_2;
  DataMuxIn5(14) <= intdelay_out_15_2;
  DataMuxIn5(15) <= intdelay_out_16_2;

  intdelay_1_3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        intdelay_1_reg_48 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_49 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_50 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_51 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_52 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_53 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_54 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_55 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_56 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_57 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_58 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_59 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_60 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_61 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_62 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_63 <= (OTHERS => to_unsigned(16#00#, 8));
      ELSIF enb = '1' AND padShift = '1' THEN
        intdelay_1_reg_48(0) <= intdelay_out_1_2;
        intdelay_1_reg_48(1) <= intdelay_1_reg_48(0);
        intdelay_1_reg_49(0) <= intdelay_out_2_2;
        intdelay_1_reg_49(1) <= intdelay_1_reg_49(0);
        intdelay_1_reg_50(0) <= intdelay_out_3_2;
        intdelay_1_reg_50(1) <= intdelay_1_reg_50(0);
        intdelay_1_reg_51(0) <= intdelay_out_4_2;
        intdelay_1_reg_51(1) <= intdelay_1_reg_51(0);
        intdelay_1_reg_52(0) <= intdelay_out_5_2;
        intdelay_1_reg_52(1) <= intdelay_1_reg_52(0);
        intdelay_1_reg_53(0) <= intdelay_out_6_2;
        intdelay_1_reg_53(1) <= intdelay_1_reg_53(0);
        intdelay_1_reg_54(0) <= intdelay_out_7_2;
        intdelay_1_reg_54(1) <= intdelay_1_reg_54(0);
        intdelay_1_reg_55(0) <= intdelay_out_8_2;
        intdelay_1_reg_55(1) <= intdelay_1_reg_55(0);
        intdelay_1_reg_56(0) <= intdelay_out_9_2;
        intdelay_1_reg_56(1) <= intdelay_1_reg_56(0);
        intdelay_1_reg_57(0) <= intdelay_out_10_2;
        intdelay_1_reg_57(1) <= intdelay_1_reg_57(0);
        intdelay_1_reg_58(0) <= intdelay_out_11_2;
        intdelay_1_reg_58(1) <= intdelay_1_reg_58(0);
        intdelay_1_reg_59(0) <= intdelay_out_12_2;
        intdelay_1_reg_59(1) <= intdelay_1_reg_59(0);
        intdelay_1_reg_60(0) <= intdelay_out_13_2;
        intdelay_1_reg_60(1) <= intdelay_1_reg_60(0);
        intdelay_1_reg_61(0) <= intdelay_out_14_2;
        intdelay_1_reg_61(1) <= intdelay_1_reg_61(0);
        intdelay_1_reg_62(0) <= intdelay_out_15_2;
        intdelay_1_reg_62(1) <= intdelay_1_reg_62(0);
        intdelay_1_reg_63(0) <= intdelay_out_16_2;
        intdelay_1_reg_63(1) <= intdelay_1_reg_63(0);
      END IF;
    END IF;
  END PROCESS intdelay_1_3_process;

  intdelay_out_1_3 <= intdelay_1_reg_48(1);
  intdelay_out_2_3 <= intdelay_1_reg_49(1);
  intdelay_out_3_3 <= intdelay_1_reg_50(1);
  intdelay_out_4_3 <= intdelay_1_reg_51(1);
  intdelay_out_5_3 <= intdelay_1_reg_52(1);
  intdelay_out_6_3 <= intdelay_1_reg_53(1);
  intdelay_out_7_3 <= intdelay_1_reg_54(1);
  intdelay_out_8_3 <= intdelay_1_reg_55(1);
  intdelay_out_9_3 <= intdelay_1_reg_56(1);
  intdelay_out_10_3 <= intdelay_1_reg_57(1);
  intdelay_out_11_3 <= intdelay_1_reg_58(1);
  intdelay_out_12_3 <= intdelay_1_reg_59(1);
  intdelay_out_13_3 <= intdelay_1_reg_60(1);
  intdelay_out_14_3 <= intdelay_1_reg_61(1);
  intdelay_out_15_3 <= intdelay_1_reg_62(1);
  intdelay_out_16_3 <= intdelay_1_reg_63(1);

  DataMuxIn6(0) <= intdelay_out_1_3;
  DataMuxIn6(1) <= intdelay_out_2_3;
  DataMuxIn6(2) <= intdelay_out_3_3;
  DataMuxIn6(3) <= intdelay_out_4_3;
  DataMuxIn6(4) <= intdelay_out_5_3;
  DataMuxIn6(5) <= intdelay_out_6_3;
  DataMuxIn6(6) <= intdelay_out_7_3;
  DataMuxIn6(7) <= intdelay_out_8_3;
  DataMuxIn6(8) <= intdelay_out_9_3;
  DataMuxIn6(9) <= intdelay_out_10_3;
  DataMuxIn6(10) <= intdelay_out_11_3;
  DataMuxIn6(11) <= intdelay_out_12_3;
  DataMuxIn6(12) <= intdelay_out_13_3;
  DataMuxIn6(13) <= intdelay_out_14_3;
  DataMuxIn6(14) <= intdelay_out_15_3;
  DataMuxIn6(15) <= intdelay_out_16_3;

  intdelay_1_4_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        intdelay_1_reg_64 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_65 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_66 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_67 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_68 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_69 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_70 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_71 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_72 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_73 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_74 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_75 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_76 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_77 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_78 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_79 <= (OTHERS => to_unsigned(16#00#, 8));
      ELSIF enb = '1' AND padShift = '1' THEN
        intdelay_1_reg_64(0) <= intdelay_out_1_3;
        intdelay_1_reg_64(1) <= intdelay_1_reg_64(0);
        intdelay_1_reg_65(0) <= intdelay_out_2_3;
        intdelay_1_reg_65(1) <= intdelay_1_reg_65(0);
        intdelay_1_reg_66(0) <= intdelay_out_3_3;
        intdelay_1_reg_66(1) <= intdelay_1_reg_66(0);
        intdelay_1_reg_67(0) <= intdelay_out_4_3;
        intdelay_1_reg_67(1) <= intdelay_1_reg_67(0);
        intdelay_1_reg_68(0) <= intdelay_out_5_3;
        intdelay_1_reg_68(1) <= intdelay_1_reg_68(0);
        intdelay_1_reg_69(0) <= intdelay_out_6_3;
        intdelay_1_reg_69(1) <= intdelay_1_reg_69(0);
        intdelay_1_reg_70(0) <= intdelay_out_7_3;
        intdelay_1_reg_70(1) <= intdelay_1_reg_70(0);
        intdelay_1_reg_71(0) <= intdelay_out_8_3;
        intdelay_1_reg_71(1) <= intdelay_1_reg_71(0);
        intdelay_1_reg_72(0) <= intdelay_out_9_3;
        intdelay_1_reg_72(1) <= intdelay_1_reg_72(0);
        intdelay_1_reg_73(0) <= intdelay_out_10_3;
        intdelay_1_reg_73(1) <= intdelay_1_reg_73(0);
        intdelay_1_reg_74(0) <= intdelay_out_11_3;
        intdelay_1_reg_74(1) <= intdelay_1_reg_74(0);
        intdelay_1_reg_75(0) <= intdelay_out_12_3;
        intdelay_1_reg_75(1) <= intdelay_1_reg_75(0);
        intdelay_1_reg_76(0) <= intdelay_out_13_3;
        intdelay_1_reg_76(1) <= intdelay_1_reg_76(0);
        intdelay_1_reg_77(0) <= intdelay_out_14_3;
        intdelay_1_reg_77(1) <= intdelay_1_reg_77(0);
        intdelay_1_reg_78(0) <= intdelay_out_15_3;
        intdelay_1_reg_78(1) <= intdelay_1_reg_78(0);
        intdelay_1_reg_79(0) <= intdelay_out_16_3;
        intdelay_1_reg_79(1) <= intdelay_1_reg_79(0);
      END IF;
    END IF;
  END PROCESS intdelay_1_4_process;

  intdelay_out_1_4 <= intdelay_1_reg_64(1);
  intdelay_out_2_4 <= intdelay_1_reg_65(1);
  intdelay_out_3_4 <= intdelay_1_reg_66(1);
  intdelay_out_4_4 <= intdelay_1_reg_67(1);
  intdelay_out_5_4 <= intdelay_1_reg_68(1);
  intdelay_out_6_4 <= intdelay_1_reg_69(1);
  intdelay_out_7_4 <= intdelay_1_reg_70(1);
  intdelay_out_8_4 <= intdelay_1_reg_71(1);
  intdelay_out_9_4 <= intdelay_1_reg_72(1);
  intdelay_out_10_4 <= intdelay_1_reg_73(1);
  intdelay_out_11_4 <= intdelay_1_reg_74(1);
  intdelay_out_12_4 <= intdelay_1_reg_75(1);
  intdelay_out_13_4 <= intdelay_1_reg_76(1);
  intdelay_out_14_4 <= intdelay_1_reg_77(1);
  intdelay_out_15_4 <= intdelay_1_reg_78(1);
  intdelay_out_16_4 <= intdelay_1_reg_79(1);

  DataMuxIn7(0) <= intdelay_out_1_4;
  DataMuxIn7(1) <= intdelay_out_2_4;
  DataMuxIn7(2) <= intdelay_out_3_4;
  DataMuxIn7(3) <= intdelay_out_4_4;
  DataMuxIn7(4) <= intdelay_out_5_4;
  DataMuxIn7(5) <= intdelay_out_6_4;
  DataMuxIn7(6) <= intdelay_out_7_4;
  DataMuxIn7(7) <= intdelay_out_8_4;
  DataMuxIn7(8) <= intdelay_out_9_4;
  DataMuxIn7(9) <= intdelay_out_10_4;
  DataMuxIn7(10) <= intdelay_out_11_4;
  DataMuxIn7(11) <= intdelay_out_12_4;
  DataMuxIn7(12) <= intdelay_out_13_4;
  DataMuxIn7(13) <= intdelay_out_14_4;
  DataMuxIn7(14) <= intdelay_out_15_4;
  DataMuxIn7(15) <= intdelay_out_16_4;

  intdelay_1_5_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        intdelay_1_reg_80 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_81 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_82 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_83 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_84 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_85 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_86 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_87 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_88 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_89 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_90 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_91 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_92 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_93 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_94 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_95 <= (OTHERS => to_unsigned(16#00#, 8));
      ELSIF enb = '1' AND padShift = '1' THEN
        intdelay_1_reg_80(0) <= intdelay_out_1_4;
        intdelay_1_reg_80(1) <= intdelay_1_reg_80(0);
        intdelay_1_reg_81(0) <= intdelay_out_2_4;
        intdelay_1_reg_81(1) <= intdelay_1_reg_81(0);
        intdelay_1_reg_82(0) <= intdelay_out_3_4;
        intdelay_1_reg_82(1) <= intdelay_1_reg_82(0);
        intdelay_1_reg_83(0) <= intdelay_out_4_4;
        intdelay_1_reg_83(1) <= intdelay_1_reg_83(0);
        intdelay_1_reg_84(0) <= intdelay_out_5_4;
        intdelay_1_reg_84(1) <= intdelay_1_reg_84(0);
        intdelay_1_reg_85(0) <= intdelay_out_6_4;
        intdelay_1_reg_85(1) <= intdelay_1_reg_85(0);
        intdelay_1_reg_86(0) <= intdelay_out_7_4;
        intdelay_1_reg_86(1) <= intdelay_1_reg_86(0);
        intdelay_1_reg_87(0) <= intdelay_out_8_4;
        intdelay_1_reg_87(1) <= intdelay_1_reg_87(0);
        intdelay_1_reg_88(0) <= intdelay_out_9_4;
        intdelay_1_reg_88(1) <= intdelay_1_reg_88(0);
        intdelay_1_reg_89(0) <= intdelay_out_10_4;
        intdelay_1_reg_89(1) <= intdelay_1_reg_89(0);
        intdelay_1_reg_90(0) <= intdelay_out_11_4;
        intdelay_1_reg_90(1) <= intdelay_1_reg_90(0);
        intdelay_1_reg_91(0) <= intdelay_out_12_4;
        intdelay_1_reg_91(1) <= intdelay_1_reg_91(0);
        intdelay_1_reg_92(0) <= intdelay_out_13_4;
        intdelay_1_reg_92(1) <= intdelay_1_reg_92(0);
        intdelay_1_reg_93(0) <= intdelay_out_14_4;
        intdelay_1_reg_93(1) <= intdelay_1_reg_93(0);
        intdelay_1_reg_94(0) <= intdelay_out_15_4;
        intdelay_1_reg_94(1) <= intdelay_1_reg_94(0);
        intdelay_1_reg_95(0) <= intdelay_out_16_4;
        intdelay_1_reg_95(1) <= intdelay_1_reg_95(0);
      END IF;
    END IF;
  END PROCESS intdelay_1_5_process;

  intdelay_out_1_5 <= intdelay_1_reg_80(1);
  intdelay_out_2_5 <= intdelay_1_reg_81(1);
  intdelay_out_3_5 <= intdelay_1_reg_82(1);
  intdelay_out_4_5 <= intdelay_1_reg_83(1);
  intdelay_out_5_5 <= intdelay_1_reg_84(1);
  intdelay_out_6_5 <= intdelay_1_reg_85(1);
  intdelay_out_7_5 <= intdelay_1_reg_86(1);
  intdelay_out_8_5 <= intdelay_1_reg_87(1);
  intdelay_out_9_5 <= intdelay_1_reg_88(1);
  intdelay_out_10_5 <= intdelay_1_reg_89(1);
  intdelay_out_11_5 <= intdelay_1_reg_90(1);
  intdelay_out_12_5 <= intdelay_1_reg_91(1);
  intdelay_out_13_5 <= intdelay_1_reg_92(1);
  intdelay_out_14_5 <= intdelay_1_reg_93(1);
  intdelay_out_15_5 <= intdelay_1_reg_94(1);
  intdelay_out_16_5 <= intdelay_1_reg_95(1);

  DataMuxIn8(0) <= intdelay_out_1_5;
  DataMuxIn8(1) <= intdelay_out_2_5;
  DataMuxIn8(2) <= intdelay_out_3_5;
  DataMuxIn8(3) <= intdelay_out_4_5;
  DataMuxIn8(4) <= intdelay_out_5_5;
  DataMuxIn8(5) <= intdelay_out_6_5;
  DataMuxIn8(6) <= intdelay_out_7_5;
  DataMuxIn8(7) <= intdelay_out_8_5;
  DataMuxIn8(8) <= intdelay_out_9_5;
  DataMuxIn8(9) <= intdelay_out_10_5;
  DataMuxIn8(10) <= intdelay_out_11_5;
  DataMuxIn8(11) <= intdelay_out_12_5;
  DataMuxIn8(12) <= intdelay_out_13_5;
  DataMuxIn8(13) <= intdelay_out_14_5;
  DataMuxIn8(14) <= intdelay_out_15_5;
  DataMuxIn8(15) <= intdelay_out_16_5;

  intdelay_1_6_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset = '1' THEN
        intdelay_1_reg_96 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_97 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_98 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_99 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_100 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_101 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_102 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_103 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_104 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_105 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_106 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_107 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_108 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_109 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_110 <= (OTHERS => to_unsigned(16#00#, 8));
        intdelay_1_reg_111 <= (OTHERS => to_unsigned(16#00#, 8));
      ELSIF enb = '1' AND padShift = '1' THEN
        intdelay_1_reg_96(0) <= intdelay_out_1_5;
        intdelay_1_reg_96(1) <= intdelay_1_reg_96(0);
        intdelay_1_reg_97(0) <= intdelay_out_2_5;
        intdelay_1_reg_97(1) <= intdelay_1_reg_97(0);
        intdelay_1_reg_98(0) <= intdelay_out_3_5;
        intdelay_1_reg_98(1) <= intdelay_1_reg_98(0);
        intdelay_1_reg_99(0) <= intdelay_out_4_5;
        intdelay_1_reg_99(1) <= intdelay_1_reg_99(0);
        intdelay_1_reg_100(0) <= intdelay_out_5_5;
        intdelay_1_reg_100(1) <= intdelay_1_reg_100(0);
        intdelay_1_reg_101(0) <= intdelay_out_6_5;
        intdelay_1_reg_101(1) <= intdelay_1_reg_101(0);
        intdelay_1_reg_102(0) <= intdelay_out_7_5;
        intdelay_1_reg_102(1) <= intdelay_1_reg_102(0);
        intdelay_1_reg_103(0) <= intdelay_out_8_5;
        intdelay_1_reg_103(1) <= intdelay_1_reg_103(0);
        intdelay_1_reg_104(0) <= intdelay_out_9_5;
        intdelay_1_reg_104(1) <= intdelay_1_reg_104(0);
        intdelay_1_reg_105(0) <= intdelay_out_10_5;
        intdelay_1_reg_105(1) <= intdelay_1_reg_105(0);
        intdelay_1_reg_106(0) <= intdelay_out_11_5;
        intdelay_1_reg_106(1) <= intdelay_1_reg_106(0);
        intdelay_1_reg_107(0) <= intdelay_out_12_5;
        intdelay_1_reg_107(1) <= intdelay_1_reg_107(0);
        intdelay_1_reg_108(0) <= intdelay_out_13_5;
        intdelay_1_reg_108(1) <= intdelay_1_reg_108(0);
        intdelay_1_reg_109(0) <= intdelay_out_14_5;
        intdelay_1_reg_109(1) <= intdelay_1_reg_109(0);
        intdelay_1_reg_110(0) <= intdelay_out_15_5;
        intdelay_1_reg_110(1) <= intdelay_1_reg_110(0);
        intdelay_1_reg_111(0) <= intdelay_out_16_5;
        intdelay_1_reg_111(1) <= intdelay_1_reg_111(0);
      END IF;
    END IF;
  END PROCESS intdelay_1_6_process;

  intdelay_out_1_6 <= intdelay_1_reg_96(1);
  intdelay_out_2_6 <= intdelay_1_reg_97(1);
  intdelay_out_3_6 <= intdelay_1_reg_98(1);
  intdelay_out_4_6 <= intdelay_1_reg_99(1);
  intdelay_out_5_6 <= intdelay_1_reg_100(1);
  intdelay_out_6_6 <= intdelay_1_reg_101(1);
  intdelay_out_7_6 <= intdelay_1_reg_102(1);
  intdelay_out_8_6 <= intdelay_1_reg_103(1);
  intdelay_out_9_6 <= intdelay_1_reg_104(1);
  intdelay_out_10_6 <= intdelay_1_reg_105(1);
  intdelay_out_11_6 <= intdelay_1_reg_106(1);
  intdelay_out_12_6 <= intdelay_1_reg_107(1);
  intdelay_out_13_6 <= intdelay_1_reg_108(1);
  intdelay_out_14_6 <= intdelay_1_reg_109(1);
  intdelay_out_15_6 <= intdelay_1_reg_110(1);
  intdelay_out_16_6 <= intdelay_1_reg_111(1);

  DataMuxIn9(0) <= intdelay_out_1_6;
  DataMuxIn9(1) <= intdelay_out_2_6;
  DataMuxIn9(2) <= intdelay_out_3_6;
  DataMuxIn9(3) <= intdelay_out_4_6;
  DataMuxIn9(4) <= intdelay_out_5_6;
  DataMuxIn9(5) <= intdelay_out_6_6;
  DataMuxIn9(6) <= intdelay_out_7_6;
  DataMuxIn9(7) <= intdelay_out_8_6;
  DataMuxIn9(8) <= intdelay_out_9_6;
  DataMuxIn9(9) <= intdelay_out_10_6;
  DataMuxIn9(10) <= intdelay_out_11_6;
  DataMuxIn9(11) <= intdelay_out_12_6;
  DataMuxIn9(12) <= intdelay_out_13_6;
  DataMuxIn9(13) <= intdelay_out_14_6;
  DataMuxIn9(14) <= intdelay_out_15_6;
  DataMuxIn9(15) <= intdelay_out_16_6;

  mux_output : PROCESS (DataMuxIn1, DataMuxIn1_16, DataMuxIn2, DataMuxIn3, DataMuxIn4, DataMuxIn5,
       DataMuxIn6, DataMuxIn7, DataMuxIn8, DataMuxIn9, horPadCount_unsigned)
  BEGIN
    IF horPadCount_unsigned = to_unsigned(16#000#, 11) THEN 
      dataVector_tmp <= DataMuxIn1;
    ELSIF horPadCount_unsigned = to_unsigned(16#001#, 11) THEN 
      dataVector_tmp <= DataMuxIn1_16;
    ELSIF horPadCount_unsigned = to_unsigned(16#002#, 11) THEN 
      dataVector_tmp <= DataMuxIn2;
    ELSIF horPadCount_unsigned = to_unsigned(16#003#, 11) THEN 
      dataVector_tmp <= DataMuxIn3;
    ELSIF horPadCount_unsigned = to_unsigned(16#004#, 11) THEN 
      dataVector_tmp <= DataMuxIn4;
    ELSIF horPadCount_unsigned = to_unsigned(16#005#, 11) THEN 
      dataVector_tmp <= DataMuxIn5;
    ELSIF horPadCount_unsigned = to_unsigned(16#006#, 11) THEN 
      dataVector_tmp <= DataMuxIn6;
    ELSIF horPadCount_unsigned = to_unsigned(16#007#, 11) THEN 
      dataVector_tmp <= DataMuxIn7;
    ELSIF horPadCount_unsigned = to_unsigned(16#008#, 11) THEN 
      dataVector_tmp <= DataMuxIn8;
    ELSE 
      dataVector_tmp <= DataMuxIn9;
    END IF;
  END PROCESS mux_output;


  outputgen: FOR k IN 0 TO 15 GENERATE
    dataVector(k) <= std_logic_vector(dataVector_tmp(k));
  END GENERATE;

END rtl;

